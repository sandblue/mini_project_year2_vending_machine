library verilog;
use verilog.vl_types.all;
entity eightBitToBcd_vlg_vec_tst is
end eightBitToBcd_vlg_vec_tst;
