library verilog;
use verilog.vl_types.all;
entity MuxTwo_vlg_vec_tst is
end MuxTwo_vlg_vec_tst;
