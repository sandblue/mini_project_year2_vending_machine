library verilog;
use verilog.vl_types.all;
entity debounce_switch_vlg_vec_tst is
end debounce_switch_vlg_vec_tst;
