library ieee;
use ieee.std_logic_1164.all;

entity detectRisingEdge is
    port(input)