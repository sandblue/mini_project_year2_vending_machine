library verilog;
use verilog.vl_types.all;
entity divid_clk_vlg_vec_tst is
end divid_clk_vlg_vec_tst;
