library verilog;
use verilog.vl_types.all;
entity debounce_switch_vlg_check_tst is
    port(
        result          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end debounce_switch_vlg_check_tst;
