library verilog;
use verilog.vl_types.all;
entity vending_mach_vlg_vec_tst is
end vending_mach_vlg_vec_tst;
