library verilog;
use verilog.vl_types.all;
entity process_price_vlg_vec_tst is
end process_price_vlg_vec_tst;
