library verilog;
use verilog.vl_types.all;
entity calValue_vlg_vec_tst is
end calValue_vlg_vec_tst;
