library verilog;
use verilog.vl_types.all;
entity insertComplete_vlg_check_tst is
    port(
        output_buzzer_on: in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end insertComplete_vlg_check_tst;
