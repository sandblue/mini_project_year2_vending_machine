library verilog;
use verilog.vl_types.all;
entity open_buzzer_vlg_vec_tst is
end open_buzzer_vlg_vec_tst;
