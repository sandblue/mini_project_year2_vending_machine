library verilog;
use verilog.vl_types.all;
entity insertComplete_vlg_vec_tst is
end insertComplete_vlg_vec_tst;
