library verilog;
use verilog.vl_types.all;
entity insertCoin_vlg_vec_tst is
end insertCoin_vlg_vec_tst;
