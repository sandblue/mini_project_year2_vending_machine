library verilog;
use verilog.vl_types.all;
entity detectRisingEdge_vlg_vec_tst is
end detectRisingEdge_vlg_vec_tst;
