library verilog;
use verilog.vl_types.all;
entity clk_to_selecter_vlg_vec_tst is
end clk_to_selecter_vlg_vec_tst;
