library verilog;
use verilog.vl_types.all;
entity clk_to_selecter_vlg_check_tst is
    port(
        o               : in     vl_logic;
        ob              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end clk_to_selecter_vlg_check_tst;
