library verilog;
use verilog.vl_types.all;
entity open_buzzer_vlg_check_tst is
    port(
        out_buzzer      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end open_buzzer_vlg_check_tst;
