library verilog;
use verilog.vl_types.all;
entity detectRisingEdge_vlg_check_tst is
    port(
        o               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end detectRisingEdge_vlg_check_tst;
