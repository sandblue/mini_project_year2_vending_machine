library verilog;
use verilog.vl_types.all;
entity divid_clk_vlg_check_tst is
    port(
        clk_after       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end divid_clk_vlg_check_tst;
