library verilog;
use verilog.vl_types.all;
entity buyMode_vlg_check_tst is
    port(
        mode            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end buyMode_vlg_check_tst;
