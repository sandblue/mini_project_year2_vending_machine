library verilog;
use verilog.vl_types.all;
entity buyMode_vlg_vec_tst is
end buyMode_vlg_vec_tst;
